
----------------------------------------------------------------------------------
-- MIT License
-- 
-- Copyright (c) 2022 Martin Skriver
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
----------------------------------------------------------------------------------
-- Company: University of Southern Denmark
-- Engineer: Martin Skriver
-- Contact: maskr@mmmi.sdu.dk maskr09@gmail.com
--
-- Description: 
-- Memory inst for positive signal for HEIST
--
----------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------
-- Libraries 
-----------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VComponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

-----------------------------------------------------------------------------------------------------
-- Ports and generics
-----------------------------------------------------------------------------------------------------
entity pos_sig_bram_mem_interface is
    Port ( clk_in           : in STD_LOGIC;
           addr_in          : in STD_LOGIC_VECTOR (11 downto 0);
           data_out         : out STD_LOGIC_VECTOR (7 downto 0));
end pos_sig_bram_mem_interface;

architecture Behavioral of pos_sig_bram_mem_interface is

begin
BRAM_TDP_MACRO_inst : BRAM_TDP_MACRO
    generic map (
        BRAM_SIZE           => "36Kb",        -- Target BRAM, "18Kb" or "36Kb"
        DEVICE              => "7SERIES",       -- Target Device: "VIRTEX5", "VIRTEX6", "7SERIES", "SPARTAN6"
        DOA_REG             => 0,               -- Optional port A output register (0 or 1)
        DOB_REG             => 0,               -- Optional port B output register (0 or 1)
        INIT_A              => X"000000000",    -- Initial values on A output port
        INIT_B              => X"000000000",    -- Initial values on B output port
        INIT_FILE           => "NONE",
        READ_WIDTH_A        => 8,    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH_B        => 8,    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY",
        -- "GENERATE_X_ONLY" or "NONE"
        SRVAL_A             => X"000000000",    -- Set/Reset value for A port output
        SRVAL_B             => X"000000000",    -- Set/Reset value for B port output
        WRITE_MODE_A        => "WRITE_FIRST",   -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        WRITE_MODE_B        => "WRITE_FIRST",   -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        WRITE_WIDTH_A       => 8,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        WRITE_WIDTH_B       => 8,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")

--      Burst level:  resolution check
--      Last adress:  0b000000100000

        -- The following INIT_xx declarations specify the initial contents of the RAM
        INIT_00 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFAAFFFF00FF80FFC0FFE0FFF0FFF8FFFCFFFEFF",
        INIT_01 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000", 
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",

        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INIT_xx are valid when configured as 36Kb
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INITP_xx are for the parity bits
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INIT_xx are valid when configured as 36Kb
        INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
    )

----      Burst level:  2.0
----      Last adress:  0b111110100000

--        -- The following INIT_xx declarations specify the initial contents of the RAM
--        INIT_00 => X"c03ff03ff801ff00ff803fe01ff007f803ff01ff801f803ff83f8001f83ffffc",
--        INIT_01 => X"ff803fc01ff00ff803ff01ff801f803ff83f8003f83ffffcaac3ffff3ffe07ff",
--        INIT_02 => X"01ff01ffc01f803ff83fc001f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_03 => X"f83fc001f83ffffeaac0ffff1fff07ffe01ff01ffc01ff00ff801fe01ff007f8",
--        INIT_04 => X"aac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_05 => X"e01ff01ff801ff00ff803fe01ff007f803ff01ffc01f803ff83fc001f83ffffc",
--        INIT_06 => X"ffc01fe01ff807f801ff00ffc00fc03ffc3fc001f83ffffeaac0ffff3fff07ff",
--        INIT_07 => X"01ff01ffc00fc03ff83fc001f83ffffcaae07fff1fff03ffe01ff00ffc01ff00", 
--        INIT_08 => X"f83f8003f83ffffcaac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f8",
--        INIT_09 => X"aac0fffe3ffe07ffc03ff01ff803fe01ff803fc03ff00ff003ff01ff801f803f",
--        INIT_0A => X"e01ff80ffc01ff00ffc01fe01ff807f801ff00ffc00fc03ffc3fc001f83ffffe",
--        INIT_0B => X"ff803fc03ff00ff003ff01ff801f803ff83f8003f87ffffcaae07fff1fff03ff",
--        INIT_0C => X"03ff01ffc01f803ff83fc001f83ffffcaac0fffe3ffe07ffc03ff01ff803fe01",
--        INIT_0D => X"f83fc001f83ffffcaac07fff1fff07ffe01ff01ffc01ff00ff801fe01ff007f8",
--        INIT_0E => X"aac0ffff1fff07ffe01ff01ffc01ff00ff801fe01ff007f803ff01ffc01f803f",
--        INIT_0F => X"e01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03ffc3fc001f83ffffe",
--        INIT_10 => X"ff803fe01ff007f803ff01ff801f803ff83f8001f83ffffcaae07fff1fff03ff",
--        INIT_11 => X"01ff00ffc00fc03ffc3fc001f83ffffeaac0ffff3ffe07ffc03ff01ff801fe00",
--        INIT_12 => X"f83fc001f83ffffeaae07fff1fff03ffe01ff00ffc01ff00ffc01fe01ff807f8",
--        INIT_13 => X"aac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_14 => X"e01ff00ffc01ff00ffc01fe01ff807f801ff01ffc00f803ff83fc001f83ffffc",
--        INIT_15 => X"ff803fc01ff00ff803ff01ff801f803ff83f8001f83ffffcaac07fff1fff07ff",
--        INIT_16 => X"03ff01ffc01f803ff83fc001f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_17 => X"fc3fc001f83ffffeaac0ffff1fff07ffe01ff01ff801ff00ff803fe01ff007f8",
--        INIT_18 => X"aac07fff1fff03ffe01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_19 => X"e01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03ffc3fc001f83ffffe",
--        INIT_1A => X"ff801fe01ff007f803ff01ffc01f803ff83fc001f83ffffcaae07fff1fff03ff",

--        INIT_1B => X"03ff01ff801f803ff83f8001f83ffffcaac07fff1fff07ffe01ff01ffc01ff00",
--        INIT_1C => X"f83fc001f83ffffcaac0ffff3ffe07ffc03ff01ff801fe00ff803fe01ff007f8",
--        INIT_1D => X"aac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_1E => X"c03ff01ff801fe00ff803fe01ff007f803ff01ff801f803ff83f8001f83ffffc",
--        INIT_1F => X"ff803fc01ff00ff003ff01ff801f803ff83f8001f83ffffcaac0ffff3ffe07ff",
--        INIT_20 => X"01ff00ffc00fc03ff83fc001f83ffffeaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_21 => X"f83fc001f83ffffcaac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f8",
--        INIT_22 => X"aac0ffff1fff07ffe01ff01ff801ff00ff803fe01ff007f803ff01ffc01f803f",
--        INIT_23 => X"e01ff01ff801ff00ff801fe01ff007f803ff01ffc01f803ff83fc001f83ffffc",
--        INIT_24 => X"ff803fe01ff007f803ff01ff801f803ff83f8001f83ffffcaac07fff1fff07ff",
--        INIT_25 => X"01ff00ffc00fc03ffc3fc001f83ffffeaac0ffff3ffe07ffc03ff01ff801fe00",
--        INIT_26 => X"f83fc001f83ffffcaae07fff1fff03ffe01ff00ffc01ff00ffc01fe01ff807f8",
--        INIT_27 => X"aac07fff1fff07ffe01ff01ffc01ff00ff801fe01ff007f801ff01ffc01f803f",
--        INIT_28 => X"c03ff01ff803fe01ff803fc03ff00ff003ff01ff801f803ff83f8003f83ffffc",
--        INIT_29 => X"ffc01fe01ff807f801ff01ffc00fc03ff83fc001f83ffffcaac0fffe3ffe07ff",
--        INIT_2A => X"03ff01ff801f803ff83f8001f83ffffcaac07fff1fff07ffe01ff01ffc01ff00",
--        INIT_2B => X"fc3fc001f83ffffeaac0ffff3fff07ffe01ff01ff801ff00ff803fe01ff007f8",
--        INIT_2C => X"aac07fff1fff03ffe01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_2D => X"e01ff01ffc01ff00ff801fe01ff007f801ff01ffc01f803ff83fc001f83ffffc",
--        INIT_2E => X"ff803fe01ff007f803ff01ff801f803ff83fc001f83ffffcaac07fff1fff07ff",
--        INIT_2F => X"01ff01ffc01f803ff83fc001f83ffffcaac0ffff1fff07ffe01ff01ff801ff00",
--        INIT_30 => X"f83f8001f83ffffcaac07fff1fff07ffe01ff01ff801ff00ff801fe01ff007f8",
--        INIT_31 => X"aac0ffff3ffe07ffc03ff01ff801fe00ff803fe01ff007f803ff01ff801f803f",
--        INIT_32 => X"e01ff01ffc01ff00ff801fe01ff007f801ff01ffc01f803ff83fc001f83ffffc",
--        INIT_33 => X"ff803fc03ff00ff003ff01ff801f803ff83f8003f83ffffcaac0ffff1fff07ff",
--        INIT_34 => X"03ff01ff801f803ff83f8003f87ffffcaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_35 => X"f83f8003f83ffffcaac0fffe3ffe07ffc03ff01ff803fe01ff803fc03ff00ff0",
--        INIT_36 => X"aac0fffe3ffe07ffc03ff01ff801fe01ff803fc03ff00ff003ff01ff801f803f",
--        INIT_37 => X"c03ff01ff801fe00ff803fc01ff007f803ff01ff801f803ff83f8001f83ffffc",
--        INIT_38 => X"ff803fe01ff007f803ff01ff801f803ff83f8001f83ffffcaac0ffff3ffe07ff",
--        INIT_39 => X"03ff01ffc01f803ff83fc001f83ffffcaac0ffff3fff07ffe01ff01ff801ff00",
--        INIT_3A => X"fc3fc001f83ffffeaac0ffff1fff07ffe01ff01ff801ff00ff803fe01ff007f8",
--        INIT_3B => X"aae07fff1fff03ffe01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_3C => X"e01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03ffc3fc001f83ffffe",
--        INIT_3D => X"ff803fc03ff00ff003ff01ff801f803ff83f8003f83ffffcaae07fff1fff03ff",
--        INIT_3E => X"03ff01ffc01f803ff83fc001f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_3F => X"f83f8003f87ffffcaac0ffff1fff07ffe01ff01ffc01ff00ff801fe01ff007f8",
--        -- The next set of INIT_xx are valid when configured as 36Kb
--        INIT_40 => X"aac0fffe3ffe07ffc03ff01ff803fe01ff803fc03ff00ff003fe01ff801f807f",
--        INIT_41 => X"e01ff01ff801ff00ff803fe01ff007f803ff01ffc01f803ff83fc001f83ffffc",
--        INIT_42 => X"ff803fe01ff007f803ff01ffc01f803ff83fc001f83ffffcaac0ffff1fff07ff",
--        INIT_43 => X"01ff00ffc00fc03ff83fc001f83ffffeaac0ffff1fff07ffe01ff01ff801ff00",
--        INIT_44 => X"f83fc001f83ffffcaac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f8",
--        INIT_45 => X"aac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f801ff01ffc00f803f",
--        INIT_46 => X"e01ff01ff801ff00ffc01fe01ff007f801ff01ffc01f803ff83fc001f83ffffc",
--        INIT_47 => X"ffc01fe01ff807f801ff01ffc00f803ff83fc001f83ffffcaac0ffff1fff07ff",
--        INIT_48 => X"03ff01ff801f803ff83f8003f83ffffcaac07fff1fff07ffe01ff00ffc01ff00",
--        INIT_49 => X"f83f8003f83ffffcaac0fffe3ffe07ffc03ff01ff803fe01ff803fc03ff00ff0",
--        INIT_4A => X"aac0fffe3ffe07ffc03ff01ff803fe01ff803fc03ff00ff003ff01ff801f803f",
--        INIT_4B => X"c03ff01ff801fe00ff803fe01ff007f803ff01ff801f803ff83f8001f83ffffc",
--        INIT_4C => X"ff803fc01ff007f003ff01ff801f803ff83f8001f83ffffcaac0ffff3ffe07ff",
--        INIT_4D => X"03ff01ff801f803ff83f8001f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_4E => X"fc3fc001f83ffffeaac0ffff3fff07ffe01ff01ff801ff00ff803fe01ff007f8",
--        INIT_4F => X"aae07fff1fff03ffe01ff80ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_50 => X"e01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03ffc3fc001f83ffffe",
--        INIT_51 => X"ff803fe01ff007f803ff01ffc01f803ff83fc001f83ffffcaae07fff1fff03ff",
--        INIT_52 => X"03ff01ff801f803ff83f8003f83ffffcaac0ffff1fff07ffe01ff01ff801ff00",
--        INIT_53 => X"f83f8003f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01ff803fc03ff00ff0",
--        INIT_54 => X"aac0fffe3ffe07ffc03ff01ff801fe01ff803fc03ff00ff003ff01ff801f803f",
--        INIT_55 => X"e01ff01ff801ff00ff803fe01ff007f803ff01ffc01f803ff83fc001f83ffffc",
--        INIT_56 => X"ffc01fe01ff807f801ff80ffc00fc03ffc1fc001fc3ffffeaac0ffff1fff07ff",
--        INIT_57 => X"03ff01ff801f803ff83f8003f83ffffcaae07fff1fff03ffe01ff80ffc01ff00",
--        INIT_58 => X"f83fc001f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01ff803fc01ff00ff0",
--        INIT_59 => X"aac07fff1fff07ffe01ff01ffc01ff00ffc01fe01ff007f801ff01ffc00fc03f",
--        INIT_5A => X"c03ff01ff801fe00ff803fc01ff007f803ff01ff801f803ff83f8001f83ffffc",
--        INIT_5B => X"ff803fe01ff007f801ff01ffc01f803ff83fc001f83ffffcaac0ffff3ffe07ff",
--        INIT_5C => X"03ff01ff801f803ff83f8003f83ffffcaac07fff1fff07ffe01ff01ff801ff00",
--        INIT_5D => X"f83f8001f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01ff803fc03ff00ff0",
--        INIT_5E => X"aa83fffe7ffe0fffc07ff03ff801ff01ff803fc01ff00ff803ff01ff801f803f",
--        INIT_5F => X"c03ff01ff801fe01ff803fc01ff00ff803ff01ff801f803ff83f8001f83ffffc",
--        INIT_60 => X"ff803fe01ff007f803ff01ffc01f803ff83fc001f83ffffcaac0ffff3ffe07ff",
--        INIT_61 => X"03ff01ff801f803ff83f8003f83ffffcaac0ffff1fff07ffe01ff01ff801ff00",
--        INIT_62 => X"f83f8001f83ffffcaac0fffe3ffe07ffc03ff01ff801fe01ff803fc01ff00ff0",
--        INIT_63 => X"aac0ffff3ffe07ffc01ff01ff801fe00ff803fe01ff007f803ff01ff801f803f",
--        INIT_64 => X"c03ff01ff803fe01ff803fc03ff00ff003ff01ff801f803ff83f8003f83ffffc",
--        INIT_65 => X"ffc01fe01ff807f801ff80ffc00fc03ffc3fc001fc3ffffeaac0fffe3ffe07ff",
--        INIT_66 => X"01ff01ffc00f803ff83fc001f83ffffcaae07fff1fff03ffe01ff80ffc01ff00",
--        INIT_67 => X"f83f8001f83ffffcaac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f8",
--        INIT_68 => X"aac0ffff3ffe07ffc03ff01ff801fe00ff803fe01ff007f803ff01ff801f803f",
--        INIT_69 => X"e01ff80ffc01ff00ffc01fe01ff807f801ff80ffc00fc03ffc3fc001fc3ffffe",
--        INIT_6A => X"ff803fe01ff007f803ff01ff801f803ff83f8001f83ffffcaae07fff1fff03ff",
--        INIT_6B => X"03ff01ff801f803ff83f8003f83ffffcaac0ffff3ffe07ffc01ff01ff801ff00",
--        INIT_6C => X"fc3fc001f83ffffeaac0fffe3ffe07ffc03ff01ff801fe01ff803fc03ff00ff0",
--        INIT_6D => X"aae07fff1fff03ffe01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03f",
--        INIT_6E => X"e01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03ff83fc001f83ffffe",
--        INIT_6F => X"ff801fe01ff807f801ff01ffc01f803ff83fc001f83ffffcaac07fff1fff07ff",
--        INIT_70 => X"03ff01ff801f803ff83f8003f87ffffcaac07fff1fff07ffe01ff01ffc01ff00",
--        INIT_71 => X"f83fc001f83ffffcaac0fffe3ffe07ffc03ff01ff803fe01ff803fc03ff00ff0",
--        INIT_72 => X"aac0ffff1fff07ffe01ff01ff801ff00ff803fe01ff007f803ff01ffc01f803f",
--        INIT_73 => X"e01ff00ffc01ff00ffc01fe01ff807f801ff00ffc00fc03ffc3fc001fc3ffffe",
--        INIT_74 => X"ff803fc01ff00ff003ff01ff801f803ff83f8001f83ffffcaae07fff1fff03ff",
--        INIT_75 => X"03ff01ff801f803ff83f8003f87ffffcaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_76 => X"f83fc001f83ffffcaac0fffe3ffe07ffc03ff01ff803fe01ff803fc03ff00ff0",
--        INIT_77 => X"aac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f801ff01ffc00fc03f",
--        INIT_78 => X"c03ff01ff801fe01ff803fc01ff00ff003ff01ff801f803ff83f8001f83ffffc",
--        INIT_79 => X"ff803fc01ff007f803ff01ff801f803ff83f8001f83ffffcaac0fffe3ffe07ff",
--        INIT_7A => X"01ff00ffc00fc03ffc3fc001f83ffffeaac0fffe3ffe07ffc03ff01ff801fe01",
--        INIT_7B => X"f83fc001f83ffffcaac07fff1fff07ffe01ff00ffc01ff00ffc01fe01ff807f8",
--        INIT_7C => X"aac0ffff3fff07ffe01ff01ff801ff00ff803fe01ff007f803ff01ffc01f803f",
--        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
--        -- The next set of INITP_xx are for the parity bits
--        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        -- The next set of INIT_xx are valid when configured as 36Kb
--        INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
--    )

    port map (
        DOA => data_out,             -- Output port-A data, width defined by READ_WIDTH_A parameter
        DOB => open,             -- Output port-B data, width defined by READ_WIDTH_B parameter
        ADDRA => addr_in,         -- Input port-A address, width defined by Port A depth
        ADDRB => "000000000000",         -- Input port-B address, width defined by Port B depth
        CLKA => clk_in,           -- 1-bit input port-A clock
        CLKB => clk_in,           -- 1-bit input port-B clock
        DIA => (others => '0'),             -- Input port-A data, width defined by WRITE_WIDTH_A parameter
        DIB => (others => '0'),             -- Input port-B data, width defined by WRITE_WIDTH_B parameter
        ENA => '1',             -- 1-bit input port-A enable
        ENB => '0',             -- 1-bit input port-B enable
--        REGCEA => REGCEA_in,       -- 1-bit input port-A output register enable
--        REGCEB => REGCEB_in,       -- 1-bit input port-B output register enable
        REGCEA => '0',       -- 1-bit input port-A output register enable
        REGCEB => '0',       -- 1-bit input port-B output register enable
        RSTA => '0',           -- 1-bit input port-A reset
        RSTB => '0',           -- 1-bit input port-B reset
        WEA => "0",             -- Input port-A write enable, width defined by Port A depth
        WEB => "0"              -- Input port-B write enable, width defined by Port B depth
    );


end Behavioral;
