
----------------------------------------------------------------------------------
-- MIT License
-- 
-- Copyright (c) 2022 Martin Skriver
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.
----------------------------------------------------------------------------------
-- Company: University of Southern Denmark
-- Engineer: Martin Skriver
-- Contact: maskr@mmmi.sdu.dk maskr09@gmail.com
--
-- Description: 
-- Memory inst negative signal HEIST
--
----------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------
-- Libraries 
-----------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VComponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

-----------------------------------------------------------------------------------------------------
-- Ports and generics
-----------------------------------------------------------------------------------------------------
entity neg_sig_bram_mem_interface is
    Port ( clk_in           : in STD_LOGIC;
           addr_in          : in STD_LOGIC_VECTOR (11 downto 0);
           data_out         : out STD_LOGIC_VECTOR (7 downto 0));
end neg_sig_bram_mem_interface;

architecture Behavioral of neg_sig_bram_mem_interface is

begin
BRAM_TDP_MACRO_inst : BRAM_TDP_MACRO 
    generic map (
        BRAM_SIZE           => "36Kb",        -- Target BRAM, "18Kb" or "36Kb"
        DEVICE              => "7SERIES",       -- Target Device: "VIRTEX5", "VIRTEX6", "7SERIES", "SPARTAN6"
        DOA_REG             => 0,               -- Optional port A output register (0 or 1)
        DOB_REG             => 0,               -- Optional port B output register (0 or 1)
        INIT_A              => X"000000000",    -- Initial values on A output port
        INIT_B              => X"000000000",    -- Initial values on B output port
        INIT_FILE           => "NONE",
        READ_WIDTH_A        => 8,    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH_B        => 8,    -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY",
        -- "GENERATE_X_ONLY" or "NONE"
        SRVAL_A             => X"000000000",    -- Set/Reset value for A port output
        SRVAL_B             => X"000000000",    -- Set/Reset value for B port output
        WRITE_MODE_A        => "WRITE_FIRST",   -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        WRITE_MODE_B        => "WRITE_FIRST",   -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
        WRITE_WIDTH_A       => 8,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
        WRITE_WIDTH_B       => 8,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")


--      Burst level:  resolution check
--      Last adress:  0b000000100000

        -- The following INIT_xx declarations specify the initial contents of the RAM
        INIT_00 => X"0000000000000000000000000000AA00FF007F003F001F000F00070003000100",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000", 
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",

        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INIT_xx are valid when configured as 36Kb
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INITP_xx are for the parity bits
        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        -- The next set of INIT_xx are valid when configured as 36Kb
        INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
    )
    
----      Burst level:  2.0
----      Last adress:  0b111110010110
--        -- The following INIT_xx declarations specify the initial contents of the RAM
--        INIT_00 => X"c001e000fc001fc00ff003f801ff007f003fe01ff801f803ff83f8001f87ffe7",
--        INIT_01 => X"0fc007f801fc00ff007f801ff00ff800f803ff83fc001f83fff3aae000000007",
--        INIT_02 => X"00ff007f801ff00ffc00f801ff83fc001f83fff3aa7800000007e000f0007e00",
--        INIT_03 => X"f00ff800f803ff83fc001f83fff3aa7800000003e000f0007e000fe007f801fc",
--        INIT_04 => X"ff83fc001f83fff7aa7800000007e000f0007e000fc007f801fc00ff007f801f",
--        INIT_05 => X"fff3aa7800000007e000f0007e001fc007f801fc01ff007f801ff00ff800f803",
--        INIT_06 => X"0003e000f0007e000fe007f801fc00ff007f801ff00ffc00f801ff83fc001f83",
--        INIT_07 => X"7e000fc007f801fc00ff007f801ff00ff800f803ff83fc001f83fff3aa780000", 
--        INIT_08 => X"01fc01ff007f001ff01ff800f803ff83f8001f83ffe7aa7800000007e000f000",
--        INIT_09 => X"001ff01ff800f803ff83f8001f83ffe7aa7800000007e000f0007e001fc007f8",
--        INIT_0A => X"f803ff83f8001f87ffe7aa7800000007e000f0007e001fc007f801fc01ff007f",
--        INIT_0B => X"1f83fff3aa7000000007c001f000fe001fc00ff803fc01fe007f003fe01ff801",
--        INIT_0C => X"00000003e000f0007e000fe007f801fc00ff007f801ff00ff800f803ff83fc00",
--        INIT_0D => X"f0007e001fc007f801fc01ff007f001ff01ff800f803ff83f8001f83ffe7aa78",
--        INIT_0E => X"07f801fc00ff007f801ff00ffc00fc01ff81fc001f83fff3aa7800000007e000", 
--        INIT_0F => X"007f801ff00ffc00fc01ffc1fc001f83fff3aa7800000003e000f8007f000fe0",
--        INIT_10 => X"f800f803ff83f8001f83ffe7aa7800000003e000f8007f000fe007f801fc00ff",
--        INIT_11 => X"f8001f83ffe7aa7800000007e000f0007e001fc007f801fc01ff007f801ff01f",
--        INIT_12 => X"aa7000000007c001f000fe001fc00ff803fc01ff007f003fe01ff801f803ff83",
--        INIT_13 => X"e000f0007e000fe007f801fc00ff007f801ff00ffc00f801ff83fc001f83fff3",
--        INIT_14 => X"1fc007f801fc01ff007f001ff01ff800f803ff83f8001f83ffe7aa7800000003",
--        INIT_15 => X"01ff007f801ff00ff800f803ff83fc001f83fff7aa7800000007e000f0007e00",
--        INIT_16 => X"f01ff800f803ff83f8001f83ffe7aa7800000007e000f0007e001fc007f801fc",
--        INIT_17 => X"ff83fc001f83fff7aa7800000007e000f0007e001fc007f801fc01ff007f001f",
--        INIT_18 => X"fff7aa7800000007e000f0007e001fc007f801fc01ff007f801ff00ff800f803",
--        INIT_19 => X"0007e000f0007e001fc007f801fc01ff007f801ff00ff800f803ff83fc001f83",
--        INIT_1A => X"7e001fc00ff801fc01ff007f003ff01ff801f803ff83f8001f83ffe7aa780000",
--        INIT_1B => X"01fc01ff007f801ff01ff800f803ff83f8001f83fff7aa7000000007e001f000",
--        INIT_1C => X"003ff01ff801f803ff83f8001f83ffe7aa7800000007e000f0007e001fc007f8",
--        INIT_1D => X"f803ff83f8001f83ffe7aa7000000007e001f000fe001fc00ff801fc01ff007f",
--        INIT_1E => X"1f83ffe7aa7800000007e000f0007e001fc007f801fc01ff007f001ff01ff800",
--        INIT_1F => X"00000007e000f0007e001fc007f801fc01ff007f003ff01ff800f803ff83f800",
--        INIT_20 => X"f0007e000fe007f801fc00ff007f801ff00ff800f801ff83fc001f83fff3aa78",
--        INIT_21 => X"07f801fc01ff007f001ff01ff800f803ff83f8001f83ffe7aa7800000007e000",
--        INIT_22 => X"007f003ff01ff801f803ff83f8001f83ffe7aa7800000007e000f0007e001fc0",
--        INIT_23 => X"f800f803ff83f8001f83ffe7aa7000000007c001f000fe001fc00ff803fc01ff",
--        INIT_24 => X"f8001f83ffe7aa7800000007e000f0007e001fc007f801fc01ff007f001ff01f",
--        INIT_25 => X"aaf000000007c001f000fe001fc00ff803f801fe007f003fe01ff801f803ff83",
--        INIT_26 => X"c001f000fe001fc00ff003f801fe007f003fe01ff801f803ff83f8003f87ffe7",
--        INIT_27 => X"1fc00ff801fc01ff007f003ff01ff800f803ff83f8001f83ffe7aaf000000007",
--        INIT_28 => X"00ff007f801ff00ff800f803ff83fc001f83fff3aa7800000007e000f0007e00",
--        INIT_29 => X"f01ff801f803ff83f8001f83ffe7aa7800000007e000f0007e000fc007f801fc",
--        INIT_2A => X"ffc1fc001f83fff3aa7800000007e000f0007e001fc00ff801fc01ff007f003f",
--        INIT_2B => X"ffe7aa7800000003e000f8007e000fe007f801fc00ff007f801ff00ffc00fc01",
--        INIT_2C => X"0007c001f000fe001fc00ff803fc01ff007f003ff01ff801f803ff83f8001f83",
--        INIT_2D => X"fe001fc00ff003f801fe007f003fe01ff801f803ff83f8001f87ffe7aa700000",
--        INIT_2E => X"01fc01ff007f003ff01ff801f803ff83f8001f83ffe7aaf000000007c001f000",
--        INIT_2F => X"003fe01ff801f803ff83f8001f87ffe7aa7800000007e001f000fe001fc00ff8",
--        INIT_30 => X"f803ff83fc001f83fff3aaf000000007c001f000fe001fc00ff003f801fe007f",
--        INIT_31 => X"1f87ffe7aa7800000007e000f0007e000fe007f801fc00ff007f801ff00ff800",
--        INIT_32 => X"00000007c001f000fe001fc00ff803fc01fe007f003fe01ff801f803ff83f800",
--        INIT_33 => X"f0007e001fc00ff801fc01ff007f003ff01ff800f803ff83f8001f83ffe7aaf0",
--        INIT_34 => X"0ff801fc01ff007f003ff01ff801f803ff83f8001f83ffe7aa7800000007e000",
--        INIT_35 => X"00ff003fe01ff801f803ff83f8001f87ffe7aa7000000007e001f0007e001fc0",
--        INIT_36 => X"f800f803ff83fc001f83fff3aaf000000007c001f000fe001fc00ff003f801fe",
--        INIT_37 => X"fc001f83fff3aa7800000007e000f0007e000fc007f801fc00ff007f801ff00f",
--        INIT_38 => X"aa7800000003e000f0007e000fe007f801fc00ff007f801ff00ff800f801ff83",
--        INIT_39 => X"c001f000fe001fc00ff803fc01ff007f003fe01ff801f803ff83f8001f83ffe7",
--        INIT_3A => X"1fc007f801fc01ff007f801ff00ff800f803ff83fc001f83fff3aa7000000007",
--        INIT_3B => X"01ff007f003ff01ff801f803ff83f8001f83ffe7aa7800000007e000f0007e00",
--        INIT_3C => X"e01ff801f803ff83f8001f83ffe7aa7000000007c001f000fe001fc00ff801fc",
--        INIT_3D => X"ff83fc001f83fff7aa7000000007c001f000fe001fc00ff803fc01ff007f003f",
--        INIT_3E => X"ffe7aa7800000007e000f0007e001fc007f801fc00ff007f801ff00ff800f803",
--        INIT_3F => X"0007c001f000fe001fc00ff803fc01ff007f003fe01ff801f803ff83f8001f83",
--        -- The next set of INIT_xx are valid when configured as 36Kb
--        INIT_40 => X"7e001fc007f801fc01ff007f801ff00ff800f803ff83fc001f83fff7aa700000",
--        INIT_41 => X"01fc00ff007f801ff00ffc00f801ff83fc001f83fff3aa7800000007e000f000",
--        INIT_42 => X"801ff00ff800f801ff83fc001f83fff3aa7800000003e000f0007e000fe007f8",
--        INIT_43 => X"f803ff83f8001f83ffe7aa7800000007e000f0007e000fe007f801fc00ff007f",
--        INIT_44 => X"1f83fff7aa7000000007e001f000fe001fc00ff801fc01ff007f003ff01ff801",
--        INIT_45 => X"00000007e000f0007e001fc007f801fc01ff007f801ff00ff800f803ff83fc00",
--        INIT_46 => X"f0007e001fc007f801fc01ff007f003ff01ff800f803ff83f8001f83ffe7aa78",
--        INIT_47 => X"0ff803fc01ff007f003fe01ff801f803ff83f8001f83ffe7aa7800000007e000",
--        INIT_48 => X"007f003ff01ff800f803ff83f8001f83ffe7aa7000000007c001f000fe001fc0",
--        INIT_49 => X"f801f803ff83f8001f87ffe7aa7800000007e000f0007e001fc007f801fc01ff",
--        INIT_4A => X"fc001f83fff3aaf000000007c001f000fe001fc00ff803f801fe007f003fe01f",
--        INIT_4B => X"aa7800000003e000f0007e000fe007f801fc00ff007f801ff00ffc00fc01ff81",
--        INIT_4C => X"c001f000fc001fc00ff003f801fe00ff003fe01ff801f803ff83f8003f07ffe7",
--        INIT_4D => X"1fc007f801fc01ff007f003ff01ff800f803ff83f8001f83ffe7aaf000000007",
--        INIT_4E => X"01ff007f003ff01ff801f803ff83f8001f83ffe7aa7800000007e000f0007e00",
--        INIT_4F => X"f00ff800f803ff83fc001f83fff3aa7000000007c001f000fe001fc00ff801fc",
--        INIT_50 => X"ff83f8001f83ffe7aa7800000007e000f0007e000fc007f801fc00ff007f801f",
--        INIT_51 => X"ffe7aa7800000007e000f0007e001fc007f801fc01ff007f003ff01ff800f803",
--        INIT_52 => X"0007c001f000fe001fc00ff803f801fe007f003fe01ff801f803ff83f8001f87",
--        INIT_53 => X"fe001fc00ff803fc01ff007f003fe01ff801f803ff83f8001f83ffe7aaf00000",
--        INIT_54 => X"01fc00ff007f801ff00ff800f803ff83fc001f83fff3aa7000000007c001f000",
--        INIT_55 => X"801ff00ffc00f801ff83fc001f83fff3aa7800000003e000f0007e000fe007f8",
--        INIT_56 => X"fc01ffc1fc001f83fff3aa7800000003e000f0007e000fe007f801fc00ff007f",
--        INIT_57 => X"1f83fff3aa7800000003e000f0007e000fe007f801fc00ff007f801ff00ffc00",
--        INIT_58 => X"00000007e000f0007e001fc007f801fc00ff007f801ff00ff800f803ff83fc00",
--        INIT_59 => X"f0007c001fc007f801fc01ff007f003ff01ff800f803ff83f8001f83ffe7aa78",
--        INIT_5A => X"07f801fc00ff007f801ff00ff800f803ff83fc001f83fff3aae000000007c000",
--        INIT_5B => X"007f001ff01ff800f803ff83f8001f83ffe7aa7800000007e000f0007e000fc0",
--        INIT_5C => X"fc00fc01ff81fc001f83fff3aa7800000007e000f0007e001fc007f801fc01ff",
--        INIT_5D => X"f8001f83ffe7aa7800000003e000f8007f000fe007f801fc00ff007f801ff00f",
--        INIT_5E => X"aa7800000007e000f0007e001fc007f801fc01ff007f801ff01ff800f803ff83",
--        INIT_5F => X"e000f0007e001fc007f801fc01ff007f003ff01ff800f803ff83f8001f83ffe7",
--        INIT_60 => X"1fc007f801fc01ff007f003ff01ff800f803ff83f8001f83ffe7aa7800000007",
--        INIT_61 => X"01fe007f003fe01ff801f803ff83f8001f87ffe7aa7800000007e000f0007e00",
--        INIT_62 => X"f01ff800f803ff83f8001f83ffe7aaf000000007c001f000fe001fc00ff003f8",
--        INIT_63 => X"ff83f8001f83ffe7aa7800000007e000f0007e001fc007f801fc01ff007f801f",
--        INIT_64 => X"fff7aa7000000007e000f0007e001fc007f801fc01ff007f003ff01ff800f803",
--        INIT_65 => X"0007e000f0007e001fc007f801fc01ff007f801ff00ff800f803ff83fc001f83",
--        INIT_66 => X"fe001fc00ff803fc01ff007f003fe01ff801f803ff83f8001f83ffe7aa780000",
--        INIT_67 => X"01fc00ff007f801ff00ff800f803ff83fc001f83fff7aa7000000007c001f000",
--        INIT_68 => X"801ff00ff800f803ff83fc001f83fff7aa7800000007e000f0007e001fc007f8",
--        INIT_69 => X"f803ff83f8001f83ffe7aa7800000007e000f0007e001fc007f801fc01ff007f",
--        INIT_6A => X"1f83fff3aa7800000007e000f0007e001fc007f801fc01ff007f001ff01ff800",
--        INIT_6B => X"00000003e000f0007e000fe007f801fc00ff007f801ff00ff800f801ff83fc00",
--        INIT_6C => X"f0007e000fe007f801fc00ff007f801ff00ffc00fc01ff81fc001f83fff3aa78",
--        INIT_6D => X"0ff801fc01ff007f003ff01ff801f803ff83f8001f83ffe7aa7800000003e000",
--        INIT_6E => X"007f003fe01ff801f803ff83f8001f83ffe7aa7000000007e000f0007e001fc0",
--        INIT_6F => X"f801f803ff83f8001f83ffe7aa7000000007c001f000fe001fc00ff803fc01ff",
--        INIT_70 => X"f8001f83ffe7aa7000000007c001f000fe001fc00ff803fc01ff007f003fe01f",
--        INIT_71 => X"aa7800000007e000f0007e001fc007f801fc01ff007f003ff01ff800f803ff83",
--        INIT_72 => X"e000f0007e001fc007f801fc01ff007f003ff01ff800f803ff83f8001f83ffe7",
--        INIT_73 => X"1fc00ff801fc01ff007f003ff01ff801f803ff83f8001f83ffe7aa7800000007",
--        INIT_74 => X"00ff007f801ff00ff800f801ff83fc001f83fff3aa7800000007e000f0007e00",
--        INIT_75 => X"f01ff800f803ff83f8001f83ffe7aa7800000007e000f0007e000fc007f801fc",
--        INIT_76 => X"ff83f8001f87ffe7aa7800000007e000f0007e001fc007f801fc01ff007f001f",
--        INIT_77 => X"fff3aaf000000007c001f000fe001fc00ff003f801fe007f003fe01ff801f803",
--        INIT_78 => X"0007e000f0007e000fc007f801fc00ff007f801ff00ff800f803ff83fc001f83",
--        INIT_79 => X"7e000fe007f801fc00ff007f801ff00ffc00fc01ff81fc001f83fff3aa780000",
--        INIT_7A => X"01fc01ff007f001ff00ff800f803ff83f8001f83ffe7aa7800000003e000f800",
--        INIT_7B => X"801ff00ff800f801ff83fc001f83fff3aa7800000007e000f0007e001fc007f8",
--        INIT_7C => X"00000000000000000000aa7800000003e000f0007e000fe007f801fc00ff007f",
--        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
--        -- The next set of INITP_xx are for the parity bits
--        INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        -- The next set of INIT_xx are valid when configured as 36Kb
--        INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
--        INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
--    )        
    port map (
        DOA => data_out,             -- Output port-A data, width defined by READ_WIDTH_A parameter
        DOB => open,             -- Output port-B data, width defined by READ_WIDTH_B parameter
        ADDRA => addr_in,         -- Input port-A address, width defined by Port A depth
        ADDRB => "000000000000",         -- Input port-B address, width defined by Port B depth
        CLKA => clk_in,           -- 1-bit input port-A clock
        CLKB => clk_in,           -- 1-bit input port-B clock
        DIA => (others => '0'),             -- Input port-A data, width defined by WRITE_WIDTH_A parameter
        DIB => (others => '0'),             -- Input port-B data, width defined by WRITE_WIDTH_B parameter
        ENA => '1',             -- 1-bit input port-A enable
        ENB => '0',             -- 1-bit input port-B enable
--        REGCEA => REGCEA_in,       -- 1-bit input port-A output register enable
--        REGCEB => REGCEB_in,       -- 1-bit input port-B output register enable
        REGCEA => '0',       -- 1-bit input port-A output register enable
        REGCEB => '0',       -- 1-bit input port-B output register enable
        RSTA => '0',           -- 1-bit input port-A reset
        RSTB => '0',           -- 1-bit input port-B reset
        WEA => "0",             -- Input port-A write enable, width defined by Port A depth
        WEB => "0"              -- Input port-B write enable, width defined by Port B depth
    );


end Behavioral;
